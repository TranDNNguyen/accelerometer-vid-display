module scaling();

endmodule
