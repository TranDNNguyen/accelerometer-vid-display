module top_tb();

top UUT();

endmodule
